//////////////////////////////////////////////////////////////////////////////////
// Create Date:    15:14:11 03/15/2018 
// PWM transmitter + LSK demodulator code. (RS232 serial communication with PC)
// Created by JCH
//	Pin assignment for DSP-PLUS II board (company : Libertron)
//  <Port name>		<FPGA Board name>
//		i_Clock			(internal clock)			
//		PWM_OUT				
//		PWM_ENABLE			
//		LSK_IN				
//		o_Tx_Serial			
//		o_Tx_Serial_Test
//	
// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@		FOR TAPE5		     @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@	   OPTION7 is MODIFIED @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
//
//////////////////////////////////////////////////////////////////////////////////
module LSK_v1(i_Clock,DIP_SW,LED_OUT,PWM_OUT, PWM_ENABLE, LSK_IN, o_Tx_Serial, o_Tx_Serial_Test 
    //,data_tx
	 );

	input i_Clock; 			//FPGA internal Clock = 100MHz
	input [7:0] DIP_SW;		//FPGA DIP_switch
									//DIP_SW[0] -> PWM data stream mode, 
									//DIP_SW[1:7] -> Option[0:6]
	input LSK_IN;				//Data input from LSK Module
	wire [31:0] rDATA;		//Restored DATA from LSK_rDATA function
	wire Update;				//rDATA Update signal from LSK_rDATA function
	wire [2:0] trigger_state; 			//FSM states of LSK_rDATA function
	reg  [2:0] max_trigger_state = 0;//max_trigger_state store
	
	output [7:0] LED_OUT;	//FPGA LED On/Off
	output reg PWM_OUT;		//PWM DATA stream out
	output reg PWM_ENABLE;	//Power Amp enable signal
	
	reg i_Tx_DV = 0;				//UART Enable
	reg [7:0] i_Tx_Byte = 0; 	//UART Transmit 8-bit data
	wire o_Tx_Active;				//UART active signal
	wire o_Tx_Done;				//UART finish signal
	output o_Tx_Serial;			//UART serial output,, FPGA pin(UART0_TXD) : L24
	output o_Tx_Serial_Test;	//o_Tx_Serial output test pin
	reg uart_start = 0;			//uart start signal. 'High' when rDATA[31:0] update
	reg [31:0] data_tx = 0;		//uart tx data. from rDATA[31:0]
	reg [4:0] addr_index =0;	//data_tx's address 
	
	reg [0:639] PWM_STREAM_BUFF = 1;			//PWM data stream buffer
	reg [9:0] i_Clock_count=0;
	reg [21:0] PWM_CLK_COUNT=0;
	reg PWM_CAP_END = 0;							//PWM capacitor tuning end flag
	reg PWM_CLK = 1;
	reg CLK_MAX_LED = 0;					//LED On and Off , when PWM_CLK_COUNT == PWM_CLK_COUNT_MAX
	
	//PWM data option
	wire [0:19] Option7;
	wire [0:19] Option6;
	wire [0:19] Option5;
	wire [0:19] Option4;
	wire [0:19] Option3;
	wire [0:19] Option2;
	wire [0:19] Option1;
	wire [0:19] Option0;
	
	parameter CLKS_PER_BIT = 869;
	// UART
	// Example: 10 MHz i_Clock, 115200 baud UART
	// (10000000)/(115200) = 87
	//if 100MHz clock, 115200 -> 869
	//i_Clock is internal clock in FPGA (Default : 100MHz, port # : H17)
	
	parameter [7:0] PWM_CLK_CODE = 84;										//PWM_CLK(period) = i_Clock(=10ns) * PWL_CLK_CODE // PWM_CLK_CODE >= 4	
	parameter PWM_CAP_COUNT = 0;												//MAX7060 internal capacitor tuning code. Range : 4.5pF + 0~7.75pF (0.25pF step, 32 levels)
	parameter PWM_CLK_COUNT_MAX = 22'b01_1111_1111_1111_1111_1111;	//PWM_CLK_COUNT max value
	
	parameter PWM_DATA_HIGH = 20'b0000_0000_0000_1111_1111;	//Duty 40%
	parameter PWM_DATA_LOW  = 20'b0000_0000_0000_0000_0001;	//Duty  5%
	
	//stream data(order : left to right) 
	//-> Header(16 bits) : 0110_1110_1111_0100, Data(8 bits) : Option<7:0> defaults : 0000_1110
	//Option<7> is not used in Tape2 Chip. 
	//Option<7> is used in Tape5 Chip. (For current level change)
	
	//assign Option7 = PWM_DATA_HIGH;	//default 0, no used (Tape2)
	assign Option7 = DIP_SW[1] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 0 : CURRENT_SENSOR UNIT I increase
	assign Option6 = DIP_SW[7] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 0 : IOP_RES_TOGGLE
	assign Option5 = DIP_SW[6] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 0 : LED_ON				
	assign Option4 = DIP_SW[5] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 0 : TIME<1>			
 	assign Option3 = DIP_SW[4] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 1 : TIME<0>	
	assign Option2 = DIP_SW[3] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 1 : DDS_SEL<2>
	assign Option1 = DIP_SW[2] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 1 : DDS_SEL<1>
	//assign Option0 = DIP_SW[1] ? PWM_DATA_HIGH : PWM_DATA_LOW;	//default 0 : DDS_SEL<0>
	assign Option0 = PWM_DATA_LOW;	//default 0 in Tape5
	
	assign LED_OUT[7:4] = 0;			//not used
	assign LED_OUT[0] = CLK_MAX_LED;
	assign LED_OUT[3:1] = DIP_SW[0] ? 3'b000 : max_trigger_state;	//Modeified in Tape5
	
	assign o_Tx_Serial_Test = o_Tx_Serial;	//test pin
	
	LSK_rDATA uut (
		.i_Clock(i_Clock), 
		.LSK_IN(LSK_IN), 
		.rDATA(rDATA), 
		.Update(Update),
		.trigger_state(trigger_state)
	);
		
	uart_tx my_uart_RS232(
		  .i_Clock(i_Clock),
		  .i_Tx_DV(i_Tx_DV),
		  .i_Tx_Byte(i_Tx_Byte), 
		  .o_Tx_Active(o_Tx_Active), 
		  .o_Tx_Serial(o_Tx_Serial), 
		  .o_Tx_Done(o_Tx_Done),
		  .CLKS_PER_BIT(CLKS_PER_BIT)
		  );
		
	always @(posedge i_Clock) begin
		//test code
		if(trigger_state > max_trigger_state)	max_trigger_state <= trigger_state;

		//PWM_CLK Generation
		if(i_Clock_count == PWM_CLK_CODE[7:1] - 1) begin
			PWM_CLK <= ~PWM_CLK;
			i_Clock_count <= 0;
		end
		else begin
			i_Clock_count <= i_Clock_count + 1;
		end
		
		//UART
		if(Update) begin		//rDATA[31:0] Update signal. 'High' during 1 clock cycle in LSK_rDATA function. (SAMPLE_CLK = i_Clock / 4, 25MHz)
				uart_start <= 1'b1;
				data_tx[31:0] <= rDATA[31:0];
		end
		else begin	//Update == 0
			if(uart_start) begin
				if(o_Tx_Done) begin		//o_Tx_Done 'High' when UART finishes during 1 i_Clock cycle
					i_Tx_DV <= 1'b0;
					if(addr_index < 24)	begin
						addr_index <= addr_index + 8;
					end
					else begin
						addr_index <= 0;
						uart_start <= 0;		//UART ends
					end
				end
				else begin	//o_Tx_Done == 0
					i_Tx_DV <= 1'b1;	//UART enable
					i_Tx_Byte[0] <= data_tx[31 - addr_index];		//Due to JAVA decoding code,
					i_Tx_Byte[1] <= data_tx[30 - addr_index];		//do not follow conventional UART data stream order
					i_Tx_Byte[2] <= data_tx[29 - addr_index];		//conventional : start(1-bit) - D[0:7] - stop(1-bit)
					i_Tx_Byte[3] <= data_tx[28 - addr_index];		//changed  		: start(1-bit) - D[7:0] - stop(1-bit)
					i_Tx_Byte[4] <= data_tx[27 - addr_index];
					i_Tx_Byte[5] <= data_tx[26 - addr_index];
					i_Tx_Byte[6] <= data_tx[25 - addr_index];
					i_Tx_Byte[7] <= data_tx[24 - addr_index];
				end				
			end
			else begin 	//uart_start == 0
				addr_index <= 0;
			end
		end
	end	
	
	//PWM_OUT signal generation
	always @(posedge PWM_CLK) begin
		if(DIP_SW[0] == 1'b0) begin
			PWM_ENABLE <= 1'b1;			
			PWM_CLK_COUNT <= 0;
			PWM_CAP_END <= 0;
			
			if(PWM_ENABLE == 1) PWM_OUT <= 1'b1; 
			else PWM_OUT <= 1'b0;
			
			//Data stream insertion
			PWM_STREAM_BUFF[0		:19]	<=PWM_DATA_HIGH; 		//buffer
			PWM_STREAM_BUFF[20	:39]	<=PWM_DATA_HIGH; 		
			PWM_STREAM_BUFF[40	:59]	<=PWM_DATA_HIGH; 		
			PWM_STREAM_BUFF[60	:79]	<=PWM_DATA_HIGH; 		//buffer
			PWM_STREAM_BUFF[80	:99]	<=PWM_DATA_LOW;		//Header starts
			PWM_STREAM_BUFF[100	:119]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[120	:139]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[140	:159]	<=PWM_DATA_LOW;		
			PWM_STREAM_BUFF[160	:179]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[180	:199]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[200	:219]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[220	:239]	<=PWM_DATA_LOW;		
			PWM_STREAM_BUFF[240	:259]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[260	:279]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[280	:299]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[300	:319]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[320	:339]	<=PWM_DATA_LOW;		
			PWM_STREAM_BUFF[340	:359]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[360	:379]	<=PWM_DATA_LOW;		
			PWM_STREAM_BUFF[380	:399]	<=PWM_DATA_LOW;		//Header ends
			PWM_STREAM_BUFF[400	:419]	<=Option7;				//Option<7:0> starts
			PWM_STREAM_BUFF[420	:439]	<=Option6;		
			PWM_STREAM_BUFF[440	:459]	<=Option5;		
			PWM_STREAM_BUFF[460	:479]	<=Option4;		
			PWM_STREAM_BUFF[480	:499]	<=Option3;		
			PWM_STREAM_BUFF[500	:519]	<=Option2;		
			PWM_STREAM_BUFF[520	:539]	<=Option1;		
			PWM_STREAM_BUFF[540	:559]	<=Option0;				//Option<7:0> ends 
			PWM_STREAM_BUFF[560	:579]	<=PWM_DATA_HIGH;		//buffer
			PWM_STREAM_BUFF[580	:599]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[600	:619]	<=PWM_DATA_HIGH;		
			PWM_STREAM_BUFF[620	:639]	<=PWM_DATA_HIGH;		//buffer
		end
		else begin			//DIP_SW[0] == 1 -> PWM_Mode
				if(PWM_CLK_COUNT < PWM_CLK_COUNT_MAX) begin
					PWM_CLK_COUNT <= PWM_CLK_COUNT + 1;
				end
				else begin
					PWM_CLK_COUNT <= 500;					//500 -> Àû´çÇÑ °ª
					CLK_MAX_LED <= ~CLK_MAX_LED;			//LED ON and OFF
				end
				
				//capacitor tuning code starts
				if(PWM_CLK_COUNT == 0) PWM_OUT <= 0;
				if(PWM_CLK_COUNT == 1) PWM_ENABLE <= 0;
				if(PWM_ENABLE == 0) begin
					if(PWM_CLK_COUNT-2 < 2*(PWM_CAP_COUNT+1)) begin		//PWM_CLK_COUNT-2 -> PWM_CLK_COUNT=2 starts,  
						if(PWM_OUT == 0) PWM_OUT <= 1;			 			//PWM_CAP_COUNT+1 -> first edge to reset capcitor setting value, 
						else PWM_OUT <= 0;										// 				*2 -> PWM_OUT 'H' and 'L'																					
					end
					else begin
						PWM_ENABLE <= 1;		//Enable 'H' before PWM_OUT = 'H'
						PWM_CAP_END <= 1;		//Cap tuning end flag.
					end
				end
			
				if(PWM_CAP_END && PWM_ENABLE) begin
					PWM_OUT <= 1;
					PWM_CAP_END <= 0;
				end
				//capacitor tuning code ends
				
				if(PWM_CLK_COUNT > 500) begin				//500 -> Àû´çÇÑ °ª.
					PWM_OUT <= PWM_STREAM_BUFF[0];
					PWM_STREAM_BUFF[0]  	<= PWM_STREAM_BUFF[1];		
					PWM_STREAM_BUFF[1]	<= PWM_STREAM_BUFF[2];		
					PWM_STREAM_BUFF[2]	<= PWM_STREAM_BUFF[3];		
					PWM_STREAM_BUFF[3]	<= PWM_STREAM_BUFF[4];		
					PWM_STREAM_BUFF[4]	<= PWM_STREAM_BUFF[5];		
					PWM_STREAM_BUFF[5]	<= PWM_STREAM_BUFF[6];		
					PWM_STREAM_BUFF[6]	<= PWM_STREAM_BUFF[7];		
					PWM_STREAM_BUFF[7]	<= PWM_STREAM_BUFF[8];		
					PWM_STREAM_BUFF[8]	<= PWM_STREAM_BUFF[9];		
					PWM_STREAM_BUFF[9]	<= PWM_STREAM_BUFF[10];		
					PWM_STREAM_BUFF[10]	<= PWM_STREAM_BUFF[11];		
					PWM_STREAM_BUFF[11]	<= PWM_STREAM_BUFF[12];		
					PWM_STREAM_BUFF[12]	<= PWM_STREAM_BUFF[13];		
					PWM_STREAM_BUFF[13]	<= PWM_STREAM_BUFF[14];		
					PWM_STREAM_BUFF[14]	<= PWM_STREAM_BUFF[15];		
					PWM_STREAM_BUFF[15]	<= PWM_STREAM_BUFF[16];		
					PWM_STREAM_BUFF[16]	<= PWM_STREAM_BUFF[17];		
					PWM_STREAM_BUFF[17]	<= PWM_STREAM_BUFF[18];		
					PWM_STREAM_BUFF[18]	<= PWM_STREAM_BUFF[19];		
					PWM_STREAM_BUFF[19]	<= PWM_STREAM_BUFF[20];		
					PWM_STREAM_BUFF[20]	<= PWM_STREAM_BUFF[21];		
					PWM_STREAM_BUFF[21]	<= PWM_STREAM_BUFF[22];		
					PWM_STREAM_BUFF[22]	<= PWM_STREAM_BUFF[23];		
					PWM_STREAM_BUFF[23]	<= PWM_STREAM_BUFF[24];		
					PWM_STREAM_BUFF[24]	<= PWM_STREAM_BUFF[25];		
					PWM_STREAM_BUFF[25]	<= PWM_STREAM_BUFF[26];		
					PWM_STREAM_BUFF[26]	<= PWM_STREAM_BUFF[27];		
					PWM_STREAM_BUFF[27]	<= PWM_STREAM_BUFF[28];		
					PWM_STREAM_BUFF[28]	<= PWM_STREAM_BUFF[29];		
					PWM_STREAM_BUFF[29]	<= PWM_STREAM_BUFF[30];		
					PWM_STREAM_BUFF[30]	<= PWM_STREAM_BUFF[31];		
					PWM_STREAM_BUFF[31]	<= PWM_STREAM_BUFF[32];		
					PWM_STREAM_BUFF[32]	<= PWM_STREAM_BUFF[33];		
					PWM_STREAM_BUFF[33]	<= PWM_STREAM_BUFF[34];		
					PWM_STREAM_BUFF[34]	<= PWM_STREAM_BUFF[35];		
					PWM_STREAM_BUFF[35]	<= PWM_STREAM_BUFF[36];		
					PWM_STREAM_BUFF[36]	<= PWM_STREAM_BUFF[37];		
					PWM_STREAM_BUFF[37]	<= PWM_STREAM_BUFF[38];		
					PWM_STREAM_BUFF[38]	<= PWM_STREAM_BUFF[39];		
					PWM_STREAM_BUFF[39]	<= PWM_STREAM_BUFF[40];		
					PWM_STREAM_BUFF[40]	<= PWM_STREAM_BUFF[41];		
					PWM_STREAM_BUFF[41]	<= PWM_STREAM_BUFF[42];		
					PWM_STREAM_BUFF[42]	<= PWM_STREAM_BUFF[43];		
					PWM_STREAM_BUFF[43]	<= PWM_STREAM_BUFF[44];		
					PWM_STREAM_BUFF[44]	<= PWM_STREAM_BUFF[45];		
					PWM_STREAM_BUFF[45]	<= PWM_STREAM_BUFF[46];		
					PWM_STREAM_BUFF[46]	<= PWM_STREAM_BUFF[47];		
					PWM_STREAM_BUFF[47]	<= PWM_STREAM_BUFF[48];		
					PWM_STREAM_BUFF[48]	<= PWM_STREAM_BUFF[49];		
					PWM_STREAM_BUFF[49]	<= PWM_STREAM_BUFF[50];		
					PWM_STREAM_BUFF[50]	<= PWM_STREAM_BUFF[51];		
					PWM_STREAM_BUFF[51]	<= PWM_STREAM_BUFF[52];		
					PWM_STREAM_BUFF[52]	<= PWM_STREAM_BUFF[53];		
					PWM_STREAM_BUFF[53]	<= PWM_STREAM_BUFF[54];		
					PWM_STREAM_BUFF[54]	<= PWM_STREAM_BUFF[55];		
					PWM_STREAM_BUFF[55]	<= PWM_STREAM_BUFF[56];		
					PWM_STREAM_BUFF[56]	<= PWM_STREAM_BUFF[57];		
					PWM_STREAM_BUFF[57]	<= PWM_STREAM_BUFF[58];		
					PWM_STREAM_BUFF[58]	<= PWM_STREAM_BUFF[59];		
					PWM_STREAM_BUFF[59]	<= PWM_STREAM_BUFF[60];		
					PWM_STREAM_BUFF[60]	<= PWM_STREAM_BUFF[61];		
					PWM_STREAM_BUFF[61]	<= PWM_STREAM_BUFF[62];		
					PWM_STREAM_BUFF[62]	<= PWM_STREAM_BUFF[63];		
					PWM_STREAM_BUFF[63]	<= PWM_STREAM_BUFF[64];		
					PWM_STREAM_BUFF[64]	<= PWM_STREAM_BUFF[65];		
					PWM_STREAM_BUFF[65]	<= PWM_STREAM_BUFF[66];		
					PWM_STREAM_BUFF[66]	<= PWM_STREAM_BUFF[67];		
					PWM_STREAM_BUFF[67]	<= PWM_STREAM_BUFF[68];		
					PWM_STREAM_BUFF[68]	<= PWM_STREAM_BUFF[69];		
					PWM_STREAM_BUFF[69]	<= PWM_STREAM_BUFF[70];		
					PWM_STREAM_BUFF[70]	<= PWM_STREAM_BUFF[71];		
					PWM_STREAM_BUFF[71]	<= PWM_STREAM_BUFF[72];		
					PWM_STREAM_BUFF[72]	<= PWM_STREAM_BUFF[73];		
					PWM_STREAM_BUFF[73]	<= PWM_STREAM_BUFF[74];		
					PWM_STREAM_BUFF[74]	<= PWM_STREAM_BUFF[75];		
					PWM_STREAM_BUFF[75]	<= PWM_STREAM_BUFF[76];		
					PWM_STREAM_BUFF[76]	<= PWM_STREAM_BUFF[77];		
					PWM_STREAM_BUFF[77]	<= PWM_STREAM_BUFF[78];		
					PWM_STREAM_BUFF[78]	<= PWM_STREAM_BUFF[79];		
					PWM_STREAM_BUFF[79]	<= PWM_STREAM_BUFF[80];		
					PWM_STREAM_BUFF[80]	<= PWM_STREAM_BUFF[81];		
					PWM_STREAM_BUFF[81]	<= PWM_STREAM_BUFF[82];		
					PWM_STREAM_BUFF[82]	<= PWM_STREAM_BUFF[83];		
					PWM_STREAM_BUFF[83]	<= PWM_STREAM_BUFF[84];		
					PWM_STREAM_BUFF[84]	<= PWM_STREAM_BUFF[85];		
					PWM_STREAM_BUFF[85]	<= PWM_STREAM_BUFF[86];		
					PWM_STREAM_BUFF[86]	<= PWM_STREAM_BUFF[87];		
					PWM_STREAM_BUFF[87]	<= PWM_STREAM_BUFF[88];		
					PWM_STREAM_BUFF[88]	<= PWM_STREAM_BUFF[89];		
					PWM_STREAM_BUFF[89]	<= PWM_STREAM_BUFF[90];		
					PWM_STREAM_BUFF[90]	<= PWM_STREAM_BUFF[91];		
					PWM_STREAM_BUFF[91]	<= PWM_STREAM_BUFF[92];		
					PWM_STREAM_BUFF[92]	<= PWM_STREAM_BUFF[93];		
					PWM_STREAM_BUFF[93]	<= PWM_STREAM_BUFF[94];		
					PWM_STREAM_BUFF[94]	<= PWM_STREAM_BUFF[95];		
					PWM_STREAM_BUFF[95]	<= PWM_STREAM_BUFF[96];		
					PWM_STREAM_BUFF[96]	<= PWM_STREAM_BUFF[97];		
					PWM_STREAM_BUFF[97]	<= PWM_STREAM_BUFF[98];		
					PWM_STREAM_BUFF[98]	<= PWM_STREAM_BUFF[99];		
					PWM_STREAM_BUFF[99]	<= PWM_STREAM_BUFF[100];		
					PWM_STREAM_BUFF[100]	<= PWM_STREAM_BUFF[101];		
					PWM_STREAM_BUFF[101]	<= PWM_STREAM_BUFF[102];		
					PWM_STREAM_BUFF[102]	<= PWM_STREAM_BUFF[103];		
					PWM_STREAM_BUFF[103]	<= PWM_STREAM_BUFF[104];		
					PWM_STREAM_BUFF[104]	<= PWM_STREAM_BUFF[105];		
					PWM_STREAM_BUFF[105]	<= PWM_STREAM_BUFF[106];		
					PWM_STREAM_BUFF[106]	<= PWM_STREAM_BUFF[107];		
					PWM_STREAM_BUFF[107]	<= PWM_STREAM_BUFF[108];		
					PWM_STREAM_BUFF[108]	<= PWM_STREAM_BUFF[109];		
					PWM_STREAM_BUFF[109]	<= PWM_STREAM_BUFF[110];		
					PWM_STREAM_BUFF[110]	<= PWM_STREAM_BUFF[111];		
					PWM_STREAM_BUFF[111]	<= PWM_STREAM_BUFF[112];		
					PWM_STREAM_BUFF[112]	<= PWM_STREAM_BUFF[113];		
					PWM_STREAM_BUFF[113]	<= PWM_STREAM_BUFF[114];		
					PWM_STREAM_BUFF[114]	<= PWM_STREAM_BUFF[115];		
					PWM_STREAM_BUFF[115]	<= PWM_STREAM_BUFF[116];		
					PWM_STREAM_BUFF[116]	<= PWM_STREAM_BUFF[117];		
					PWM_STREAM_BUFF[117]	<= PWM_STREAM_BUFF[118];		
					PWM_STREAM_BUFF[118]	<= PWM_STREAM_BUFF[119];		
					PWM_STREAM_BUFF[119]	<= PWM_STREAM_BUFF[120];		
					PWM_STREAM_BUFF[120]	<= PWM_STREAM_BUFF[121];		
					PWM_STREAM_BUFF[121]	<= PWM_STREAM_BUFF[122];		
					PWM_STREAM_BUFF[122]	<= PWM_STREAM_BUFF[123];		
					PWM_STREAM_BUFF[123]	<= PWM_STREAM_BUFF[124];		
					PWM_STREAM_BUFF[124]	<= PWM_STREAM_BUFF[125];		
					PWM_STREAM_BUFF[125]	<= PWM_STREAM_BUFF[126];		
					PWM_STREAM_BUFF[126]	<= PWM_STREAM_BUFF[127];		
					PWM_STREAM_BUFF[127]	<= PWM_STREAM_BUFF[128];		
					PWM_STREAM_BUFF[128]	<= PWM_STREAM_BUFF[129];		
					PWM_STREAM_BUFF[129]	<= PWM_STREAM_BUFF[130];		
					PWM_STREAM_BUFF[130]	<= PWM_STREAM_BUFF[131];		
					PWM_STREAM_BUFF[131]	<= PWM_STREAM_BUFF[132];		
					PWM_STREAM_BUFF[132]	<= PWM_STREAM_BUFF[133];		
					PWM_STREAM_BUFF[133]	<= PWM_STREAM_BUFF[134];		
					PWM_STREAM_BUFF[134]	<= PWM_STREAM_BUFF[135];		
					PWM_STREAM_BUFF[135]	<= PWM_STREAM_BUFF[136];		
					PWM_STREAM_BUFF[136]	<= PWM_STREAM_BUFF[137];		
					PWM_STREAM_BUFF[137]	<= PWM_STREAM_BUFF[138];		
					PWM_STREAM_BUFF[138]	<= PWM_STREAM_BUFF[139];		
					PWM_STREAM_BUFF[139]	<= PWM_STREAM_BUFF[140];		
					PWM_STREAM_BUFF[140]	<= PWM_STREAM_BUFF[141];		
					PWM_STREAM_BUFF[141]	<= PWM_STREAM_BUFF[142];		
					PWM_STREAM_BUFF[142]	<= PWM_STREAM_BUFF[143];		
					PWM_STREAM_BUFF[143]	<= PWM_STREAM_BUFF[144];		
					PWM_STREAM_BUFF[144]	<= PWM_STREAM_BUFF[145];		
					PWM_STREAM_BUFF[145]	<= PWM_STREAM_BUFF[146];		
					PWM_STREAM_BUFF[146]	<= PWM_STREAM_BUFF[147];		
					PWM_STREAM_BUFF[147]	<= PWM_STREAM_BUFF[148];		
					PWM_STREAM_BUFF[148]	<= PWM_STREAM_BUFF[149];		
					PWM_STREAM_BUFF[149]	<= PWM_STREAM_BUFF[150];		
					PWM_STREAM_BUFF[150]	<= PWM_STREAM_BUFF[151];		
					PWM_STREAM_BUFF[151]	<= PWM_STREAM_BUFF[152];		
					PWM_STREAM_BUFF[152]	<= PWM_STREAM_BUFF[153];		
					PWM_STREAM_BUFF[153]	<= PWM_STREAM_BUFF[154];		
					PWM_STREAM_BUFF[154]	<= PWM_STREAM_BUFF[155];		
					PWM_STREAM_BUFF[155]	<= PWM_STREAM_BUFF[156];		
					PWM_STREAM_BUFF[156]	<= PWM_STREAM_BUFF[157];		
					PWM_STREAM_BUFF[157]	<= PWM_STREAM_BUFF[158];		
					PWM_STREAM_BUFF[158]	<= PWM_STREAM_BUFF[159];		
					PWM_STREAM_BUFF[159]	<= PWM_STREAM_BUFF[160];		
					PWM_STREAM_BUFF[160]	<= PWM_STREAM_BUFF[161];		
					PWM_STREAM_BUFF[161]	<= PWM_STREAM_BUFF[162];		
					PWM_STREAM_BUFF[162]	<= PWM_STREAM_BUFF[163];		
					PWM_STREAM_BUFF[163]	<= PWM_STREAM_BUFF[164];		
					PWM_STREAM_BUFF[164]	<= PWM_STREAM_BUFF[165];		
					PWM_STREAM_BUFF[165]	<= PWM_STREAM_BUFF[166];		
					PWM_STREAM_BUFF[166]	<= PWM_STREAM_BUFF[167];		
					PWM_STREAM_BUFF[167]	<= PWM_STREAM_BUFF[168];		
					PWM_STREAM_BUFF[168]	<= PWM_STREAM_BUFF[169];		
					PWM_STREAM_BUFF[169]	<= PWM_STREAM_BUFF[170];		
					PWM_STREAM_BUFF[170]	<= PWM_STREAM_BUFF[171];		
					PWM_STREAM_BUFF[171]	<= PWM_STREAM_BUFF[172];		
					PWM_STREAM_BUFF[172]	<= PWM_STREAM_BUFF[173];		
					PWM_STREAM_BUFF[173]	<= PWM_STREAM_BUFF[174];		
					PWM_STREAM_BUFF[174]	<= PWM_STREAM_BUFF[175];		
					PWM_STREAM_BUFF[175]	<= PWM_STREAM_BUFF[176];		
					PWM_STREAM_BUFF[176]	<= PWM_STREAM_BUFF[177];		
					PWM_STREAM_BUFF[177]	<= PWM_STREAM_BUFF[178];		
					PWM_STREAM_BUFF[178]	<= PWM_STREAM_BUFF[179];		
					PWM_STREAM_BUFF[179]	<= PWM_STREAM_BUFF[180];		
					PWM_STREAM_BUFF[180]	<= PWM_STREAM_BUFF[181];		
					PWM_STREAM_BUFF[181]	<= PWM_STREAM_BUFF[182];		
					PWM_STREAM_BUFF[182]	<= PWM_STREAM_BUFF[183];		
					PWM_STREAM_BUFF[183]	<= PWM_STREAM_BUFF[184];		
					PWM_STREAM_BUFF[184]	<= PWM_STREAM_BUFF[185];		
					PWM_STREAM_BUFF[185]	<= PWM_STREAM_BUFF[186];		
					PWM_STREAM_BUFF[186]	<= PWM_STREAM_BUFF[187];		
					PWM_STREAM_BUFF[187]	<= PWM_STREAM_BUFF[188];		
					PWM_STREAM_BUFF[188]	<= PWM_STREAM_BUFF[189];		
					PWM_STREAM_BUFF[189]	<= PWM_STREAM_BUFF[190];		
					PWM_STREAM_BUFF[190]	<= PWM_STREAM_BUFF[191];		
					PWM_STREAM_BUFF[191]	<= PWM_STREAM_BUFF[192];		
					PWM_STREAM_BUFF[192]	<= PWM_STREAM_BUFF[193];		
					PWM_STREAM_BUFF[193]	<= PWM_STREAM_BUFF[194];		
					PWM_STREAM_BUFF[194]	<= PWM_STREAM_BUFF[195];		
					PWM_STREAM_BUFF[195]	<= PWM_STREAM_BUFF[196];		
					PWM_STREAM_BUFF[196]	<= PWM_STREAM_BUFF[197];		
					PWM_STREAM_BUFF[197]	<= PWM_STREAM_BUFF[198];		
					PWM_STREAM_BUFF[198]	<= PWM_STREAM_BUFF[199];		
					PWM_STREAM_BUFF[199]	<= PWM_STREAM_BUFF[200];		
					PWM_STREAM_BUFF[200]	<= PWM_STREAM_BUFF[201];		
					PWM_STREAM_BUFF[201]	<= PWM_STREAM_BUFF[202];		
					PWM_STREAM_BUFF[202]	<= PWM_STREAM_BUFF[203];		
					PWM_STREAM_BUFF[203]	<= PWM_STREAM_BUFF[204];		
					PWM_STREAM_BUFF[204]	<= PWM_STREAM_BUFF[205];		
					PWM_STREAM_BUFF[205]	<= PWM_STREAM_BUFF[206];		
					PWM_STREAM_BUFF[206]	<= PWM_STREAM_BUFF[207];		
					PWM_STREAM_BUFF[207]	<= PWM_STREAM_BUFF[208];		
					PWM_STREAM_BUFF[208]	<= PWM_STREAM_BUFF[209];		
					PWM_STREAM_BUFF[209]	<= PWM_STREAM_BUFF[210];		
					PWM_STREAM_BUFF[210]	<= PWM_STREAM_BUFF[211];		
					PWM_STREAM_BUFF[211]	<= PWM_STREAM_BUFF[212];		
					PWM_STREAM_BUFF[212]	<= PWM_STREAM_BUFF[213];		
					PWM_STREAM_BUFF[213]	<= PWM_STREAM_BUFF[214];		
					PWM_STREAM_BUFF[214]	<= PWM_STREAM_BUFF[215];		
					PWM_STREAM_BUFF[215]	<= PWM_STREAM_BUFF[216];		
					PWM_STREAM_BUFF[216]	<= PWM_STREAM_BUFF[217];		
					PWM_STREAM_BUFF[217]	<= PWM_STREAM_BUFF[218];		
					PWM_STREAM_BUFF[218]	<= PWM_STREAM_BUFF[219];		
					PWM_STREAM_BUFF[219]	<= PWM_STREAM_BUFF[220];		
					PWM_STREAM_BUFF[220]	<= PWM_STREAM_BUFF[221];		
					PWM_STREAM_BUFF[221]	<= PWM_STREAM_BUFF[222];		
					PWM_STREAM_BUFF[222]	<= PWM_STREAM_BUFF[223];		
					PWM_STREAM_BUFF[223]	<= PWM_STREAM_BUFF[224];		
					PWM_STREAM_BUFF[224]	<= PWM_STREAM_BUFF[225];		
					PWM_STREAM_BUFF[225]	<= PWM_STREAM_BUFF[226];		
					PWM_STREAM_BUFF[226]	<= PWM_STREAM_BUFF[227];		
					PWM_STREAM_BUFF[227]	<= PWM_STREAM_BUFF[228];		
					PWM_STREAM_BUFF[228]	<= PWM_STREAM_BUFF[229];		
					PWM_STREAM_BUFF[229]	<= PWM_STREAM_BUFF[230];		
					PWM_STREAM_BUFF[230]	<= PWM_STREAM_BUFF[231];		
					PWM_STREAM_BUFF[231]	<= PWM_STREAM_BUFF[232];		
					PWM_STREAM_BUFF[232]	<= PWM_STREAM_BUFF[233];		
					PWM_STREAM_BUFF[233]	<= PWM_STREAM_BUFF[234];		
					PWM_STREAM_BUFF[234]	<= PWM_STREAM_BUFF[235];		
					PWM_STREAM_BUFF[235]	<= PWM_STREAM_BUFF[236];		
					PWM_STREAM_BUFF[236]	<= PWM_STREAM_BUFF[237];		
					PWM_STREAM_BUFF[237]	<= PWM_STREAM_BUFF[238];		
					PWM_STREAM_BUFF[238]	<= PWM_STREAM_BUFF[239];		
					PWM_STREAM_BUFF[239]	<= PWM_STREAM_BUFF[240];		
					PWM_STREAM_BUFF[240]	<= PWM_STREAM_BUFF[241];		
					PWM_STREAM_BUFF[241]	<= PWM_STREAM_BUFF[242];		
					PWM_STREAM_BUFF[242]	<= PWM_STREAM_BUFF[243];		
					PWM_STREAM_BUFF[243]	<= PWM_STREAM_BUFF[244];		
					PWM_STREAM_BUFF[244]	<= PWM_STREAM_BUFF[245];		
					PWM_STREAM_BUFF[245]	<= PWM_STREAM_BUFF[246];		
					PWM_STREAM_BUFF[246]	<= PWM_STREAM_BUFF[247];		
					PWM_STREAM_BUFF[247]	<= PWM_STREAM_BUFF[248];		
					PWM_STREAM_BUFF[248]	<= PWM_STREAM_BUFF[249];		
					PWM_STREAM_BUFF[249]	<= PWM_STREAM_BUFF[250];		
					PWM_STREAM_BUFF[250]	<= PWM_STREAM_BUFF[251];		
					PWM_STREAM_BUFF[251]	<= PWM_STREAM_BUFF[252];		
					PWM_STREAM_BUFF[252]	<= PWM_STREAM_BUFF[253];		
					PWM_STREAM_BUFF[253]	<= PWM_STREAM_BUFF[254];		
					PWM_STREAM_BUFF[254]	<= PWM_STREAM_BUFF[255];		
					PWM_STREAM_BUFF[255]	<= PWM_STREAM_BUFF[256];		
					PWM_STREAM_BUFF[256]	<= PWM_STREAM_BUFF[257];		
					PWM_STREAM_BUFF[257]	<= PWM_STREAM_BUFF[258];		
					PWM_STREAM_BUFF[258]	<= PWM_STREAM_BUFF[259];		
					PWM_STREAM_BUFF[259]	<= PWM_STREAM_BUFF[260];		
					PWM_STREAM_BUFF[260]	<= PWM_STREAM_BUFF[261];		
					PWM_STREAM_BUFF[261]	<= PWM_STREAM_BUFF[262];		
					PWM_STREAM_BUFF[262]	<= PWM_STREAM_BUFF[263];		
					PWM_STREAM_BUFF[263]	<= PWM_STREAM_BUFF[264];		
					PWM_STREAM_BUFF[264]	<= PWM_STREAM_BUFF[265];		
					PWM_STREAM_BUFF[265]	<= PWM_STREAM_BUFF[266];		
					PWM_STREAM_BUFF[266]	<= PWM_STREAM_BUFF[267];		
					PWM_STREAM_BUFF[267]	<= PWM_STREAM_BUFF[268];		
					PWM_STREAM_BUFF[268]	<= PWM_STREAM_BUFF[269];		
					PWM_STREAM_BUFF[269]	<= PWM_STREAM_BUFF[270];		
					PWM_STREAM_BUFF[270]	<= PWM_STREAM_BUFF[271];		
					PWM_STREAM_BUFF[271]	<= PWM_STREAM_BUFF[272];		
					PWM_STREAM_BUFF[272]	<= PWM_STREAM_BUFF[273];		
					PWM_STREAM_BUFF[273]	<= PWM_STREAM_BUFF[274];		
					PWM_STREAM_BUFF[274]	<= PWM_STREAM_BUFF[275];		
					PWM_STREAM_BUFF[275]	<= PWM_STREAM_BUFF[276];		
					PWM_STREAM_BUFF[276]	<= PWM_STREAM_BUFF[277];		
					PWM_STREAM_BUFF[277]	<= PWM_STREAM_BUFF[278];		
					PWM_STREAM_BUFF[278]	<= PWM_STREAM_BUFF[279];		
					PWM_STREAM_BUFF[279]	<= PWM_STREAM_BUFF[280];		
					PWM_STREAM_BUFF[280]	<= PWM_STREAM_BUFF[281];		
					PWM_STREAM_BUFF[281]	<= PWM_STREAM_BUFF[282];		
					PWM_STREAM_BUFF[282]	<= PWM_STREAM_BUFF[283];		
					PWM_STREAM_BUFF[283]	<= PWM_STREAM_BUFF[284];		
					PWM_STREAM_BUFF[284]	<= PWM_STREAM_BUFF[285];		
					PWM_STREAM_BUFF[285]	<= PWM_STREAM_BUFF[286];		
					PWM_STREAM_BUFF[286]	<= PWM_STREAM_BUFF[287];		
					PWM_STREAM_BUFF[287]	<= PWM_STREAM_BUFF[288];		
					PWM_STREAM_BUFF[288]	<= PWM_STREAM_BUFF[289];		
					PWM_STREAM_BUFF[289]	<= PWM_STREAM_BUFF[290];		
					PWM_STREAM_BUFF[290]	<= PWM_STREAM_BUFF[291];		
					PWM_STREAM_BUFF[291]	<= PWM_STREAM_BUFF[292];		
					PWM_STREAM_BUFF[292]	<= PWM_STREAM_BUFF[293];		
					PWM_STREAM_BUFF[293]	<= PWM_STREAM_BUFF[294];		
					PWM_STREAM_BUFF[294]	<= PWM_STREAM_BUFF[295];		
					PWM_STREAM_BUFF[295]	<= PWM_STREAM_BUFF[296];		
					PWM_STREAM_BUFF[296]	<= PWM_STREAM_BUFF[297];		
					PWM_STREAM_BUFF[297]	<= PWM_STREAM_BUFF[298];		
					PWM_STREAM_BUFF[298]	<= PWM_STREAM_BUFF[299];		
					PWM_STREAM_BUFF[299]	<= PWM_STREAM_BUFF[300];		
					PWM_STREAM_BUFF[300]	<= PWM_STREAM_BUFF[301];		
					PWM_STREAM_BUFF[301]	<= PWM_STREAM_BUFF[302];		
					PWM_STREAM_BUFF[302]	<= PWM_STREAM_BUFF[303];		
					PWM_STREAM_BUFF[303]	<= PWM_STREAM_BUFF[304];		
					PWM_STREAM_BUFF[304]	<= PWM_STREAM_BUFF[305];		
					PWM_STREAM_BUFF[305]	<= PWM_STREAM_BUFF[306];		
					PWM_STREAM_BUFF[306]	<= PWM_STREAM_BUFF[307];		
					PWM_STREAM_BUFF[307]	<= PWM_STREAM_BUFF[308];		
					PWM_STREAM_BUFF[308]	<= PWM_STREAM_BUFF[309];		
					PWM_STREAM_BUFF[309]	<= PWM_STREAM_BUFF[310];		
					PWM_STREAM_BUFF[310]	<= PWM_STREAM_BUFF[311];		
					PWM_STREAM_BUFF[311]	<= PWM_STREAM_BUFF[312];		
					PWM_STREAM_BUFF[312]	<= PWM_STREAM_BUFF[313];		
					PWM_STREAM_BUFF[313]	<= PWM_STREAM_BUFF[314];		
					PWM_STREAM_BUFF[314]	<= PWM_STREAM_BUFF[315];		
					PWM_STREAM_BUFF[315]	<= PWM_STREAM_BUFF[316];		
					PWM_STREAM_BUFF[316]	<= PWM_STREAM_BUFF[317];		
					PWM_STREAM_BUFF[317]	<= PWM_STREAM_BUFF[318];		
					PWM_STREAM_BUFF[318]	<= PWM_STREAM_BUFF[319];		
					PWM_STREAM_BUFF[319]	<= PWM_STREAM_BUFF[320];		
					PWM_STREAM_BUFF[320]	<= PWM_STREAM_BUFF[321];		
					PWM_STREAM_BUFF[321]	<= PWM_STREAM_BUFF[322];		
					PWM_STREAM_BUFF[322]	<= PWM_STREAM_BUFF[323];		
					PWM_STREAM_BUFF[323]	<= PWM_STREAM_BUFF[324];		
					PWM_STREAM_BUFF[324]	<= PWM_STREAM_BUFF[325];		
					PWM_STREAM_BUFF[325]	<= PWM_STREAM_BUFF[326];		
					PWM_STREAM_BUFF[326]	<= PWM_STREAM_BUFF[327];		
					PWM_STREAM_BUFF[327]	<= PWM_STREAM_BUFF[328];		
					PWM_STREAM_BUFF[328]	<= PWM_STREAM_BUFF[329];		
					PWM_STREAM_BUFF[329]	<= PWM_STREAM_BUFF[330];		
					PWM_STREAM_BUFF[330]	<= PWM_STREAM_BUFF[331];		
					PWM_STREAM_BUFF[331]	<= PWM_STREAM_BUFF[332];		
					PWM_STREAM_BUFF[332]	<= PWM_STREAM_BUFF[333];		
					PWM_STREAM_BUFF[333]	<= PWM_STREAM_BUFF[334];		
					PWM_STREAM_BUFF[334]	<= PWM_STREAM_BUFF[335];		
					PWM_STREAM_BUFF[335]	<= PWM_STREAM_BUFF[336];		
					PWM_STREAM_BUFF[336]	<= PWM_STREAM_BUFF[337];		
					PWM_STREAM_BUFF[337]	<= PWM_STREAM_BUFF[338];		
					PWM_STREAM_BUFF[338]	<= PWM_STREAM_BUFF[339];		
					PWM_STREAM_BUFF[339]	<= PWM_STREAM_BUFF[340];		
					PWM_STREAM_BUFF[340]	<= PWM_STREAM_BUFF[341];		
					PWM_STREAM_BUFF[341]	<= PWM_STREAM_BUFF[342];		
					PWM_STREAM_BUFF[342]	<= PWM_STREAM_BUFF[343];		
					PWM_STREAM_BUFF[343]	<= PWM_STREAM_BUFF[344];		
					PWM_STREAM_BUFF[344]	<= PWM_STREAM_BUFF[345];		
					PWM_STREAM_BUFF[345]	<= PWM_STREAM_BUFF[346];		
					PWM_STREAM_BUFF[346]	<= PWM_STREAM_BUFF[347];		
					PWM_STREAM_BUFF[347]	<= PWM_STREAM_BUFF[348];		
					PWM_STREAM_BUFF[348]	<= PWM_STREAM_BUFF[349];		
					PWM_STREAM_BUFF[349]	<= PWM_STREAM_BUFF[350];		
					PWM_STREAM_BUFF[350]	<= PWM_STREAM_BUFF[351];		
					PWM_STREAM_BUFF[351]	<= PWM_STREAM_BUFF[352];		
					PWM_STREAM_BUFF[352]	<= PWM_STREAM_BUFF[353];		
					PWM_STREAM_BUFF[353]	<= PWM_STREAM_BUFF[354];		
					PWM_STREAM_BUFF[354]	<= PWM_STREAM_BUFF[355];		
					PWM_STREAM_BUFF[355]	<= PWM_STREAM_BUFF[356];		
					PWM_STREAM_BUFF[356]	<= PWM_STREAM_BUFF[357];		
					PWM_STREAM_BUFF[357]	<= PWM_STREAM_BUFF[358];		
					PWM_STREAM_BUFF[358]	<= PWM_STREAM_BUFF[359];		
					PWM_STREAM_BUFF[359]	<= PWM_STREAM_BUFF[360];		
					PWM_STREAM_BUFF[360]	<= PWM_STREAM_BUFF[361];		
					PWM_STREAM_BUFF[361]	<= PWM_STREAM_BUFF[362];		
					PWM_STREAM_BUFF[362]	<= PWM_STREAM_BUFF[363];		
					PWM_STREAM_BUFF[363]	<= PWM_STREAM_BUFF[364];		
					PWM_STREAM_BUFF[364]	<= PWM_STREAM_BUFF[365];		
					PWM_STREAM_BUFF[365]	<= PWM_STREAM_BUFF[366];		
					PWM_STREAM_BUFF[366]	<= PWM_STREAM_BUFF[367];		
					PWM_STREAM_BUFF[367]	<= PWM_STREAM_BUFF[368];		
					PWM_STREAM_BUFF[368]	<= PWM_STREAM_BUFF[369];		
					PWM_STREAM_BUFF[369]	<= PWM_STREAM_BUFF[370];		
					PWM_STREAM_BUFF[370]	<= PWM_STREAM_BUFF[371];		
					PWM_STREAM_BUFF[371]	<= PWM_STREAM_BUFF[372];		
					PWM_STREAM_BUFF[372]	<= PWM_STREAM_BUFF[373];		
					PWM_STREAM_BUFF[373]	<= PWM_STREAM_BUFF[374];		
					PWM_STREAM_BUFF[374]	<= PWM_STREAM_BUFF[375];		
					PWM_STREAM_BUFF[375]	<= PWM_STREAM_BUFF[376];		
					PWM_STREAM_BUFF[376]	<= PWM_STREAM_BUFF[377];		
					PWM_STREAM_BUFF[377]	<= PWM_STREAM_BUFF[378];		
					PWM_STREAM_BUFF[378]	<= PWM_STREAM_BUFF[379];		
					PWM_STREAM_BUFF[379]	<= PWM_STREAM_BUFF[380];		
					PWM_STREAM_BUFF[380]	<= PWM_STREAM_BUFF[381];		
					PWM_STREAM_BUFF[381]	<= PWM_STREAM_BUFF[382];		
					PWM_STREAM_BUFF[382]	<= PWM_STREAM_BUFF[383];		
					PWM_STREAM_BUFF[383]	<= PWM_STREAM_BUFF[384];		
					PWM_STREAM_BUFF[384]	<= PWM_STREAM_BUFF[385];		
					PWM_STREAM_BUFF[385]	<= PWM_STREAM_BUFF[386];		
					PWM_STREAM_BUFF[386]	<= PWM_STREAM_BUFF[387];		
					PWM_STREAM_BUFF[387]	<= PWM_STREAM_BUFF[388];		
					PWM_STREAM_BUFF[388]	<= PWM_STREAM_BUFF[389];		
					PWM_STREAM_BUFF[389]	<= PWM_STREAM_BUFF[390];		
					PWM_STREAM_BUFF[390]	<= PWM_STREAM_BUFF[391];		
					PWM_STREAM_BUFF[391]	<= PWM_STREAM_BUFF[392];		
					PWM_STREAM_BUFF[392]	<= PWM_STREAM_BUFF[393];		
					PWM_STREAM_BUFF[393]	<= PWM_STREAM_BUFF[394];		
					PWM_STREAM_BUFF[394]	<= PWM_STREAM_BUFF[395];		
					PWM_STREAM_BUFF[395]	<= PWM_STREAM_BUFF[396];		
					PWM_STREAM_BUFF[396]	<= PWM_STREAM_BUFF[397];		
					PWM_STREAM_BUFF[397]	<= PWM_STREAM_BUFF[398];		
					PWM_STREAM_BUFF[398]	<= PWM_STREAM_BUFF[399];		
					PWM_STREAM_BUFF[399]	<= PWM_STREAM_BUFF[400];		
					PWM_STREAM_BUFF[400]	<= PWM_STREAM_BUFF[401];		
					PWM_STREAM_BUFF[401]	<= PWM_STREAM_BUFF[402];		
					PWM_STREAM_BUFF[402]	<= PWM_STREAM_BUFF[403];		
					PWM_STREAM_BUFF[403]	<= PWM_STREAM_BUFF[404];		
					PWM_STREAM_BUFF[404]	<= PWM_STREAM_BUFF[405];		
					PWM_STREAM_BUFF[405]	<= PWM_STREAM_BUFF[406];		
					PWM_STREAM_BUFF[406]	<= PWM_STREAM_BUFF[407];		
					PWM_STREAM_BUFF[407]	<= PWM_STREAM_BUFF[408];		
					PWM_STREAM_BUFF[408]	<= PWM_STREAM_BUFF[409];		
					PWM_STREAM_BUFF[409]	<= PWM_STREAM_BUFF[410];		
					PWM_STREAM_BUFF[410]	<= PWM_STREAM_BUFF[411];		
					PWM_STREAM_BUFF[411]	<= PWM_STREAM_BUFF[412];		
					PWM_STREAM_BUFF[412]	<= PWM_STREAM_BUFF[413];		
					PWM_STREAM_BUFF[413]	<= PWM_STREAM_BUFF[414];		
					PWM_STREAM_BUFF[414]	<= PWM_STREAM_BUFF[415];		
					PWM_STREAM_BUFF[415]	<= PWM_STREAM_BUFF[416];		
					PWM_STREAM_BUFF[416]	<= PWM_STREAM_BUFF[417];		
					PWM_STREAM_BUFF[417]	<= PWM_STREAM_BUFF[418];		
					PWM_STREAM_BUFF[418]	<= PWM_STREAM_BUFF[419];		
					PWM_STREAM_BUFF[419]	<= PWM_STREAM_BUFF[420];		
					PWM_STREAM_BUFF[420]	<= PWM_STREAM_BUFF[421];		
					PWM_STREAM_BUFF[421]	<= PWM_STREAM_BUFF[422];		
					PWM_STREAM_BUFF[422]	<= PWM_STREAM_BUFF[423];		
					PWM_STREAM_BUFF[423]	<= PWM_STREAM_BUFF[424];		
					PWM_STREAM_BUFF[424]	<= PWM_STREAM_BUFF[425];		
					PWM_STREAM_BUFF[425]	<= PWM_STREAM_BUFF[426];		
					PWM_STREAM_BUFF[426]	<= PWM_STREAM_BUFF[427];		
					PWM_STREAM_BUFF[427]	<= PWM_STREAM_BUFF[428];		
					PWM_STREAM_BUFF[428]	<= PWM_STREAM_BUFF[429];		
					PWM_STREAM_BUFF[429]	<= PWM_STREAM_BUFF[430];		
					PWM_STREAM_BUFF[430]	<= PWM_STREAM_BUFF[431];		
					PWM_STREAM_BUFF[431]	<= PWM_STREAM_BUFF[432];		
					PWM_STREAM_BUFF[432]	<= PWM_STREAM_BUFF[433];		
					PWM_STREAM_BUFF[433]	<= PWM_STREAM_BUFF[434];		
					PWM_STREAM_BUFF[434]	<= PWM_STREAM_BUFF[435];		
					PWM_STREAM_BUFF[435]	<= PWM_STREAM_BUFF[436];		
					PWM_STREAM_BUFF[436]	<= PWM_STREAM_BUFF[437];		
					PWM_STREAM_BUFF[437]	<= PWM_STREAM_BUFF[438];		
					PWM_STREAM_BUFF[438]	<= PWM_STREAM_BUFF[439];		
					PWM_STREAM_BUFF[439]	<= PWM_STREAM_BUFF[440];		
					PWM_STREAM_BUFF[440]	<= PWM_STREAM_BUFF[441];		
					PWM_STREAM_BUFF[441]	<= PWM_STREAM_BUFF[442];		
					PWM_STREAM_BUFF[442]	<= PWM_STREAM_BUFF[443];		
					PWM_STREAM_BUFF[443]	<= PWM_STREAM_BUFF[444];		
					PWM_STREAM_BUFF[444]	<= PWM_STREAM_BUFF[445];		
					PWM_STREAM_BUFF[445]	<= PWM_STREAM_BUFF[446];		
					PWM_STREAM_BUFF[446]	<= PWM_STREAM_BUFF[447];		
					PWM_STREAM_BUFF[447]	<= PWM_STREAM_BUFF[448];		
					PWM_STREAM_BUFF[448]	<= PWM_STREAM_BUFF[449];		
					PWM_STREAM_BUFF[449]	<= PWM_STREAM_BUFF[450];		
					PWM_STREAM_BUFF[450]	<= PWM_STREAM_BUFF[451];		
					PWM_STREAM_BUFF[451]	<= PWM_STREAM_BUFF[452];		
					PWM_STREAM_BUFF[452]	<= PWM_STREAM_BUFF[453];		
					PWM_STREAM_BUFF[453]	<= PWM_STREAM_BUFF[454];		
					PWM_STREAM_BUFF[454]	<= PWM_STREAM_BUFF[455];		
					PWM_STREAM_BUFF[455]	<= PWM_STREAM_BUFF[456];		
					PWM_STREAM_BUFF[456]	<= PWM_STREAM_BUFF[457];		
					PWM_STREAM_BUFF[457]	<= PWM_STREAM_BUFF[458];		
					PWM_STREAM_BUFF[458]	<= PWM_STREAM_BUFF[459];		
					PWM_STREAM_BUFF[459]	<= PWM_STREAM_BUFF[460];		
					PWM_STREAM_BUFF[460]	<= PWM_STREAM_BUFF[461];		
					PWM_STREAM_BUFF[461]	<= PWM_STREAM_BUFF[462];		
					PWM_STREAM_BUFF[462]	<= PWM_STREAM_BUFF[463];		
					PWM_STREAM_BUFF[463]	<= PWM_STREAM_BUFF[464];		
					PWM_STREAM_BUFF[464]	<= PWM_STREAM_BUFF[465];		
					PWM_STREAM_BUFF[465]	<= PWM_STREAM_BUFF[466];		
					PWM_STREAM_BUFF[466]	<= PWM_STREAM_BUFF[467];		
					PWM_STREAM_BUFF[467]	<= PWM_STREAM_BUFF[468];		
					PWM_STREAM_BUFF[468]	<= PWM_STREAM_BUFF[469];		
					PWM_STREAM_BUFF[469]	<= PWM_STREAM_BUFF[470];		
					PWM_STREAM_BUFF[470]	<= PWM_STREAM_BUFF[471];		
					PWM_STREAM_BUFF[471]	<= PWM_STREAM_BUFF[472];		
					PWM_STREAM_BUFF[472]	<= PWM_STREAM_BUFF[473];		
					PWM_STREAM_BUFF[473]	<= PWM_STREAM_BUFF[474];		
					PWM_STREAM_BUFF[474]	<= PWM_STREAM_BUFF[475];		
					PWM_STREAM_BUFF[475]	<= PWM_STREAM_BUFF[476];		
					PWM_STREAM_BUFF[476]	<= PWM_STREAM_BUFF[477];		
					PWM_STREAM_BUFF[477]	<= PWM_STREAM_BUFF[478];		
					PWM_STREAM_BUFF[478]	<= PWM_STREAM_BUFF[479];		
					PWM_STREAM_BUFF[479]	<= PWM_STREAM_BUFF[480];		
					PWM_STREAM_BUFF[480]	<= PWM_STREAM_BUFF[481];		
					PWM_STREAM_BUFF[481]	<= PWM_STREAM_BUFF[482];		
					PWM_STREAM_BUFF[482]	<= PWM_STREAM_BUFF[483];		
					PWM_STREAM_BUFF[483]	<= PWM_STREAM_BUFF[484];		
					PWM_STREAM_BUFF[484]	<= PWM_STREAM_BUFF[485];		
					PWM_STREAM_BUFF[485]	<= PWM_STREAM_BUFF[486];		
					PWM_STREAM_BUFF[486]	<= PWM_STREAM_BUFF[487];		
					PWM_STREAM_BUFF[487]	<= PWM_STREAM_BUFF[488];		
					PWM_STREAM_BUFF[488]	<= PWM_STREAM_BUFF[489];		
					PWM_STREAM_BUFF[489]	<= PWM_STREAM_BUFF[490];		
					PWM_STREAM_BUFF[490]	<= PWM_STREAM_BUFF[491];		
					PWM_STREAM_BUFF[491]	<= PWM_STREAM_BUFF[492];		
					PWM_STREAM_BUFF[492]	<= PWM_STREAM_BUFF[493];		
					PWM_STREAM_BUFF[493]	<= PWM_STREAM_BUFF[494];		
					PWM_STREAM_BUFF[494]	<= PWM_STREAM_BUFF[495];		
					PWM_STREAM_BUFF[495]	<= PWM_STREAM_BUFF[496];		
					PWM_STREAM_BUFF[496]	<= PWM_STREAM_BUFF[497];		
					PWM_STREAM_BUFF[497]	<= PWM_STREAM_BUFF[498];		
					PWM_STREAM_BUFF[498]	<= PWM_STREAM_BUFF[499];		
					PWM_STREAM_BUFF[499]	<= PWM_STREAM_BUFF[500];		
					PWM_STREAM_BUFF[500]	<= PWM_STREAM_BUFF[501];		
					PWM_STREAM_BUFF[501]	<= PWM_STREAM_BUFF[502];		
					PWM_STREAM_BUFF[502]	<= PWM_STREAM_BUFF[503];		
					PWM_STREAM_BUFF[503]	<= PWM_STREAM_BUFF[504];		
					PWM_STREAM_BUFF[504]	<= PWM_STREAM_BUFF[505];		
					PWM_STREAM_BUFF[505]	<= PWM_STREAM_BUFF[506];		
					PWM_STREAM_BUFF[506]	<= PWM_STREAM_BUFF[507];		
					PWM_STREAM_BUFF[507]	<= PWM_STREAM_BUFF[508];		
					PWM_STREAM_BUFF[508]	<= PWM_STREAM_BUFF[509];		
					PWM_STREAM_BUFF[509]	<= PWM_STREAM_BUFF[510];		
					PWM_STREAM_BUFF[510]	<= PWM_STREAM_BUFF[511];		
					PWM_STREAM_BUFF[511]	<= PWM_STREAM_BUFF[512];		
					PWM_STREAM_BUFF[512]	<= PWM_STREAM_BUFF[513];		
					PWM_STREAM_BUFF[513]	<= PWM_STREAM_BUFF[514];		
					PWM_STREAM_BUFF[514]	<= PWM_STREAM_BUFF[515];		
					PWM_STREAM_BUFF[515]	<= PWM_STREAM_BUFF[516];		
					PWM_STREAM_BUFF[516]	<= PWM_STREAM_BUFF[517];		
					PWM_STREAM_BUFF[517]	<= PWM_STREAM_BUFF[518];		
					PWM_STREAM_BUFF[518]	<= PWM_STREAM_BUFF[519];		
					PWM_STREAM_BUFF[519]	<= PWM_STREAM_BUFF[520];		
					PWM_STREAM_BUFF[520]	<= PWM_STREAM_BUFF[521];		
					PWM_STREAM_BUFF[521]	<= PWM_STREAM_BUFF[522];		
					PWM_STREAM_BUFF[522]	<= PWM_STREAM_BUFF[523];		
					PWM_STREAM_BUFF[523]	<= PWM_STREAM_BUFF[524];		
					PWM_STREAM_BUFF[524]	<= PWM_STREAM_BUFF[525];		
					PWM_STREAM_BUFF[525]	<= PWM_STREAM_BUFF[526];		
					PWM_STREAM_BUFF[526]	<= PWM_STREAM_BUFF[527];		
					PWM_STREAM_BUFF[527]	<= PWM_STREAM_BUFF[528];		
					PWM_STREAM_BUFF[528]	<= PWM_STREAM_BUFF[529];		
					PWM_STREAM_BUFF[529]	<= PWM_STREAM_BUFF[530];		
					PWM_STREAM_BUFF[530]	<= PWM_STREAM_BUFF[531];		
					PWM_STREAM_BUFF[531]	<= PWM_STREAM_BUFF[532];		
					PWM_STREAM_BUFF[532]	<= PWM_STREAM_BUFF[533];		
					PWM_STREAM_BUFF[533]	<= PWM_STREAM_BUFF[534];		
					PWM_STREAM_BUFF[534]	<= PWM_STREAM_BUFF[535];		
					PWM_STREAM_BUFF[535]	<= PWM_STREAM_BUFF[536];		
					PWM_STREAM_BUFF[536]	<= PWM_STREAM_BUFF[537];		
					PWM_STREAM_BUFF[537]	<= PWM_STREAM_BUFF[538];		
					PWM_STREAM_BUFF[538]	<= PWM_STREAM_BUFF[539];		
					PWM_STREAM_BUFF[539]	<= PWM_STREAM_BUFF[540];		
					PWM_STREAM_BUFF[540]	<= PWM_STREAM_BUFF[541];		
					PWM_STREAM_BUFF[541]	<= PWM_STREAM_BUFF[542];		
					PWM_STREAM_BUFF[542]	<= PWM_STREAM_BUFF[543];		
					PWM_STREAM_BUFF[543]	<= PWM_STREAM_BUFF[544];		
					PWM_STREAM_BUFF[544]	<= PWM_STREAM_BUFF[545];		
					PWM_STREAM_BUFF[545]	<= PWM_STREAM_BUFF[546];		
					PWM_STREAM_BUFF[546]	<= PWM_STREAM_BUFF[547];		
					PWM_STREAM_BUFF[547]	<= PWM_STREAM_BUFF[548];		
					PWM_STREAM_BUFF[548]	<= PWM_STREAM_BUFF[549];		
					PWM_STREAM_BUFF[549]	<= PWM_STREAM_BUFF[550];		
					PWM_STREAM_BUFF[550]	<= PWM_STREAM_BUFF[551];		
					PWM_STREAM_BUFF[551]	<= PWM_STREAM_BUFF[552];		
					PWM_STREAM_BUFF[552]	<= PWM_STREAM_BUFF[553];		
					PWM_STREAM_BUFF[553]	<= PWM_STREAM_BUFF[554];		
					PWM_STREAM_BUFF[554]	<= PWM_STREAM_BUFF[555];		
					PWM_STREAM_BUFF[555]	<= PWM_STREAM_BUFF[556];		
					PWM_STREAM_BUFF[556]	<= PWM_STREAM_BUFF[557];		
					PWM_STREAM_BUFF[557]	<= PWM_STREAM_BUFF[558];		
					PWM_STREAM_BUFF[558]	<= PWM_STREAM_BUFF[559];		
					PWM_STREAM_BUFF[559]	<= PWM_STREAM_BUFF[560];		
					PWM_STREAM_BUFF[560]	<= PWM_STREAM_BUFF[561];		
					PWM_STREAM_BUFF[561]	<= PWM_STREAM_BUFF[562];		
					PWM_STREAM_BUFF[562]	<= PWM_STREAM_BUFF[563];		
					PWM_STREAM_BUFF[563]	<= PWM_STREAM_BUFF[564];		
					PWM_STREAM_BUFF[564]	<= PWM_STREAM_BUFF[565];		
					PWM_STREAM_BUFF[565]	<= PWM_STREAM_BUFF[566];		
					PWM_STREAM_BUFF[566]	<= PWM_STREAM_BUFF[567];		
					PWM_STREAM_BUFF[567]	<= PWM_STREAM_BUFF[568];		
					PWM_STREAM_BUFF[568]	<= PWM_STREAM_BUFF[569];		
					PWM_STREAM_BUFF[569]	<= PWM_STREAM_BUFF[570];		
					PWM_STREAM_BUFF[570]	<= PWM_STREAM_BUFF[571];		
					PWM_STREAM_BUFF[571]	<= PWM_STREAM_BUFF[572];		
					PWM_STREAM_BUFF[572]	<= PWM_STREAM_BUFF[573];		
					PWM_STREAM_BUFF[573]	<= PWM_STREAM_BUFF[574];		
					PWM_STREAM_BUFF[574]	<= PWM_STREAM_BUFF[575];		
					PWM_STREAM_BUFF[575]	<= PWM_STREAM_BUFF[576];		
					PWM_STREAM_BUFF[576]	<= PWM_STREAM_BUFF[577];		
					PWM_STREAM_BUFF[577]	<= PWM_STREAM_BUFF[578];		
					PWM_STREAM_BUFF[578]	<= PWM_STREAM_BUFF[579];		
					PWM_STREAM_BUFF[579]	<= PWM_STREAM_BUFF[580];		
					PWM_STREAM_BUFF[580]	<= PWM_STREAM_BUFF[581];		
					PWM_STREAM_BUFF[581]	<= PWM_STREAM_BUFF[582];		
					PWM_STREAM_BUFF[582]	<= PWM_STREAM_BUFF[583];		
					PWM_STREAM_BUFF[583]	<= PWM_STREAM_BUFF[584];		
					PWM_STREAM_BUFF[584]	<= PWM_STREAM_BUFF[585];		
					PWM_STREAM_BUFF[585]	<= PWM_STREAM_BUFF[586];		
					PWM_STREAM_BUFF[586]	<= PWM_STREAM_BUFF[587];		
					PWM_STREAM_BUFF[587]	<= PWM_STREAM_BUFF[588];		
					PWM_STREAM_BUFF[588]	<= PWM_STREAM_BUFF[589];		
					PWM_STREAM_BUFF[589]	<= PWM_STREAM_BUFF[590];		
					PWM_STREAM_BUFF[590]	<= PWM_STREAM_BUFF[591];		
					PWM_STREAM_BUFF[591]	<= PWM_STREAM_BUFF[592];		
					PWM_STREAM_BUFF[592]	<= PWM_STREAM_BUFF[593];		
					PWM_STREAM_BUFF[593]	<= PWM_STREAM_BUFF[594];		
					PWM_STREAM_BUFF[594]	<= PWM_STREAM_BUFF[595];		
					PWM_STREAM_BUFF[595]	<= PWM_STREAM_BUFF[596];		
					PWM_STREAM_BUFF[596]	<= PWM_STREAM_BUFF[597];		
					PWM_STREAM_BUFF[597]	<= PWM_STREAM_BUFF[598];		
					PWM_STREAM_BUFF[598]	<= PWM_STREAM_BUFF[599];		
					PWM_STREAM_BUFF[599]	<= PWM_STREAM_BUFF[600];		
					PWM_STREAM_BUFF[600]	<= PWM_STREAM_BUFF[601];		
					PWM_STREAM_BUFF[601]	<= PWM_STREAM_BUFF[602];		
					PWM_STREAM_BUFF[602]	<= PWM_STREAM_BUFF[603];		
					PWM_STREAM_BUFF[603]	<= PWM_STREAM_BUFF[604];		
					PWM_STREAM_BUFF[604]	<= PWM_STREAM_BUFF[605];		
					PWM_STREAM_BUFF[605]	<= PWM_STREAM_BUFF[606];		
					PWM_STREAM_BUFF[606]	<= PWM_STREAM_BUFF[607];		
					PWM_STREAM_BUFF[607]	<= PWM_STREAM_BUFF[608];		
					PWM_STREAM_BUFF[608]	<= PWM_STREAM_BUFF[609];		
					PWM_STREAM_BUFF[609]	<= PWM_STREAM_BUFF[610];		
					PWM_STREAM_BUFF[610]	<= PWM_STREAM_BUFF[611];		
					PWM_STREAM_BUFF[611]	<= PWM_STREAM_BUFF[612];		
					PWM_STREAM_BUFF[612]	<= PWM_STREAM_BUFF[613];		
					PWM_STREAM_BUFF[613]	<= PWM_STREAM_BUFF[614];		
					PWM_STREAM_BUFF[614]	<= PWM_STREAM_BUFF[615];		
					PWM_STREAM_BUFF[615]	<= PWM_STREAM_BUFF[616];		
					PWM_STREAM_BUFF[616]	<= PWM_STREAM_BUFF[617];		
					PWM_STREAM_BUFF[617]	<= PWM_STREAM_BUFF[618];		
					PWM_STREAM_BUFF[618]	<= PWM_STREAM_BUFF[619];		
					PWM_STREAM_BUFF[619]	<= PWM_STREAM_BUFF[620];		
					PWM_STREAM_BUFF[620]	<= PWM_STREAM_BUFF[621];		
					PWM_STREAM_BUFF[621]	<= PWM_STREAM_BUFF[622];		
					PWM_STREAM_BUFF[622]	<= PWM_STREAM_BUFF[623];		
					PWM_STREAM_BUFF[623]	<= PWM_STREAM_BUFF[624];		
					PWM_STREAM_BUFF[624]	<= PWM_STREAM_BUFF[625];		
					PWM_STREAM_BUFF[625]	<= PWM_STREAM_BUFF[626];		
					PWM_STREAM_BUFF[626]	<= PWM_STREAM_BUFF[627];		
					PWM_STREAM_BUFF[627]	<= PWM_STREAM_BUFF[628];		
					PWM_STREAM_BUFF[628]	<= PWM_STREAM_BUFF[629];		
					PWM_STREAM_BUFF[629]	<= PWM_STREAM_BUFF[630];		
					PWM_STREAM_BUFF[630]	<= PWM_STREAM_BUFF[631];		
					PWM_STREAM_BUFF[631]	<= PWM_STREAM_BUFF[632];		
					PWM_STREAM_BUFF[632]	<= PWM_STREAM_BUFF[633];		
					PWM_STREAM_BUFF[633]	<= PWM_STREAM_BUFF[634];		
					PWM_STREAM_BUFF[634]	<= PWM_STREAM_BUFF[635];		
					PWM_STREAM_BUFF[635]	<= PWM_STREAM_BUFF[636];		
					PWM_STREAM_BUFF[636]	<= PWM_STREAM_BUFF[637];		
					PWM_STREAM_BUFF[637]	<= PWM_STREAM_BUFF[638];		
					PWM_STREAM_BUFF[638]	<= PWM_STREAM_BUFF[639];		
					PWM_STREAM_BUFF[639]	<= 1;	
				end
				else begin	//PWM_CLK_COUNT <= 500
					//Data stream insertion
					PWM_STREAM_BUFF[0		:19]	<=PWM_DATA_HIGH; 		//buffer
					PWM_STREAM_BUFF[20	:39]	<=PWM_DATA_HIGH; 		
					PWM_STREAM_BUFF[40	:59]	<=PWM_DATA_HIGH; 		
					PWM_STREAM_BUFF[60	:79]	<=PWM_DATA_HIGH; 		//buffer
					PWM_STREAM_BUFF[80	:99]	<=PWM_DATA_LOW;		//Header starts
					PWM_STREAM_BUFF[100	:119]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[120	:139]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[140	:159]	<=PWM_DATA_LOW;		
					PWM_STREAM_BUFF[160	:179]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[180	:199]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[200	:219]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[220	:239]	<=PWM_DATA_LOW;		
					PWM_STREAM_BUFF[240	:259]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[260	:279]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[280	:299]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[300	:319]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[320	:339]	<=PWM_DATA_LOW;		
					PWM_STREAM_BUFF[340	:359]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[360	:379]	<=PWM_DATA_LOW;		
					PWM_STREAM_BUFF[380	:399]	<=PWM_DATA_LOW;		//Header ends
					PWM_STREAM_BUFF[400	:419]	<=Option7;				//Option<7:0> starts
					PWM_STREAM_BUFF[420	:439]	<=Option6;		
					PWM_STREAM_BUFF[440	:459]	<=Option5;		
					PWM_STREAM_BUFF[460	:479]	<=Option4;		
					PWM_STREAM_BUFF[480	:499]	<=Option3;		
					PWM_STREAM_BUFF[500	:519]	<=Option2;		
					PWM_STREAM_BUFF[520	:539]	<=Option1;		
					PWM_STREAM_BUFF[540	:559]	<=Option0;				//Option<7:0> ends 
					PWM_STREAM_BUFF[560	:579]	<=PWM_DATA_HIGH;		//buffer
					PWM_STREAM_BUFF[580	:599]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[600	:619]	<=PWM_DATA_HIGH;		
					PWM_STREAM_BUFF[620	:639]	<=PWM_DATA_HIGH;		//buffer
				end
		end
	end
endmodule
